library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity lau_block is
end lau_block;

architecture Behavioral of lau_block is

	

begin


end Behavioral;

